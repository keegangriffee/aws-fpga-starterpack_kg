`ifndef CL_PCIE_PERF
`define CL_PCIE_PERF

`define CL_NAME cl_pcie_perf

`define FPGA_LESS_RST

`endif
