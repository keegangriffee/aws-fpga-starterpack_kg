`ifndef CL_LED_DIP
`define CL_LED_DIP

`define CL_NAME cl_pcie_perf

`define FPGA_LESS_RST

`endif
